library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.functions.all;

entity char_bits is
    port(
        clk: in std_logic;
        reset: in std_logic;
        bcd: in std_logic_vector(3 downto 0);
        line_num: in std_logic_vector(width(34) - 1 downto 0);
        bitline: out std_logic_vector(0 to 25)
    );
end;

architecture behavioural of char_bits is
    type char is array(0 to 34) of std_logic_vector(0 to 25);
    
    constant zero: char := (
        "00000000001111111000000000",
        "00000000111111111110000000",
        "00000001111111111111000000",
        "00000011111111111111100000",
        "00000111111000001111110000",
        "00000111110000000111111000",
        "00001111100000000011111000",
        "00001111000000000001111100",
        "00011110000000000001111100",
        "00011110000000000000111100",
        "00011110000000000001111100",
        "00011110000000000011111110",
        "00111100000000000111111110",
        "00111100000000001111111110",
        "00111100000000111111011110",
        "00111100000001111110011110",
        "00111100000011111100011110",
        "00111100000111110000011110",
        "00111100011111100000011110",
        "00111100111111000000011110",
        "00111101111110000000011110",
        "00111111111000000000011110",
        "00111111110000000000011110",
        "00111111100000000000111110",
        "00011111000000000000111100",
        "00011110000000000000111100",
        "00011110000000000000111100",
        "00011111000000000001111000",
        "00001111100000000011111000",
        "00001111100000000111110000",
        "00000111111000001111110000",
        "00000011111111111111100000",
        "00000001111111111111000000",
        "00000000111111111110000000",
        "00000000001111111000000000");
    constant one: char := (
        "00000000000000000000000000",
        "00000000000011111000000000",
        "00000000001111111000000000",
        "00000000111111111000000000",
        "00000011111111111000000000",
        "00001111111011111000000000",
        "00011111110011111000000000",
        "00001111000011111000000000",
        "00001110000011111000000000",
        "00001000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00001111111111111111111100",
        "00001111111111111111111100",
        "00001111111111111111111100",
        "00001111111111111111111100",
        "00000000000000000000000000");
    constant two: char := (
        "00000000011111110000000000",
        "00000011111111111100000000",
        "00000111111111111110000000",
        "00001111111111111111000000",
        "00011111100000111111100000",
        "00001110000000001111100000",
        "00000100000000001111110000",
        "00000000000000000111110000",
        "00000000000000000111110000",
        "00000000000000000111110000",
        "00000000000000000111110000",
        "00000000000000000111110000",
        "00000000000000000111110000",
        "00000000000000001111110000",
        "00000000000000001111100000",
        "00000000000000001111100000",
        "00000000000000011111000000",
        "00000000000000111111000000",
        "00000000000001111110000000",
        "00000000000001111100000000",
        "00000000000011111100000000",
        "00000000000111111000000000",
        "00000000001111110000000000",
        "00000000011111100000000000",
        "00000000111111000000000000",
        "00000001111110000000000000",
        "00000011111100000000000000",
        "00000111111000000000000000",
        "00000111110000000000000000",
        "00001111100000000000000000",
        "00011111111111111111111100",
        "00011111111111111111111100",
        "00011111111111111111111100",
        "00011111111111111111111100",
        "00000000000000000000000000");
    constant three: char := (
        "00000011111111100000000000",
        "00001111111111111000000000",
        "00001111111111111110000000",
        "00001111111111111111000000",
        "00001100000000111111000000",
        "00000000000000001111100000",
        "00000000000000001111100000",
        "00000000000000000111100000",
        "00000000000000000111100000",
        "00000000000000000111100000",
        "00000000000000000111100000",
        "00000000000000000111100000",
        "00000000000000001111000000",
        "00000000000000011111000000",
        "00000000000000111110000000",
        "00000001111111111100000000",
        "00000001111111110000000000",
        "00000001111111111110000000",
        "00000001111111111111000000",
        "00000000000000011111100000",
        "00000000000000000111110000",
        "00000000000000000011111000",
        "00000000000000000001111000",
        "00000000000000000001111000",
        "00000000000000000001111000",
        "00000000000000000001111000",
        "00000000000000000001111000",
        "00000000000000000011110000",
        "00000000000000000011110000",
        "00000000000000001111110000",
        "00011000000000111111100000",
        "00011111111111111111000000",
        "00011111111111111110000000",
        "00011111111111111000000000",
        "00000111111111000000000000");
    constant four: char := (
        "00000000000000000000000000",
        "00000000000000111111000000",
        "00000000000001111111000000",
        "00000000000001111111000000",
        "00000000000011111111000000",
        "00000000000111111111000000",
        "00000000000111101111000000",
        "00000000001111101111000000",
        "00000000011111001111000000",
        "00000000011110001111000000",
        "00000000111110001111000000",
        "00000001111100001111000000",
        "00000001111000001111000000",
        "00000011111000001111000000",
        "00000111110000001111000000",
        "00000111100000001111000000",
        "00001111100000001111000000",
        "00001111000000001111000000",
        "00011110000000001111000000",
        "00111110000000001111000000",
        "00111100000000001111000000",
        "01111000000000001111000000",
        "11111000000000001111000000",
        "11111111111111111111111111",
        "11111111111111111111111111",
        "11111111111111111111111111",
        "11111111111111111111111111",
        "00000000000000001111000000",
        "00000000000000001111000000",
        "00000000000000001111000000",
        "00000000000000001111000000",
        "00000000000000001111000000",
        "00000000000000001111000000",
        "00000000000000001111000000",
        "00000000000000000000000000");
    constant five: char := (
        "00000000000000000000000000",
        "00001111111111111111100000",
        "00001111111111111111100000",
        "00001111111111111111100000",
        "00001111111111111111100000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111000000000000000000",
        "00001111111111110000000000",
        "00001111111111111100000000",
        "00001111111111111111000000",
        "00001111111111111111100000",
        "00000000000000111111110000",
        "00000000000000001111110000",
        "00000000000000000111111000",
        "00000000000000000011111000",
        "00000000000000000011111000",
        "00000000000000000011111000",
        "00000000000000000011111000",
        "00000000000000000011111000",
        "00000000000000000011111000",
        "00000000000000000111110000",
        "00000000000000001111110000",
        "00000000000000011111100000",
        "00011000000001111111000000",
        "00011111111111111110000000",
        "00011111111111111100000000",
        "00011111111111110000000000",
        "00000111111111000000000000");
    constant six: char := (
        "00000000000000000000000000",
        "00000000000000111111110000",
        "00000000000111111111110000",
        "00000000011111111111110000",
        "00000001111111111111110000",
        "00000011111111000000000000",
        "00000011111000000000000000",
        "00000111110000000000000000",
        "00001111100000000000000000",
        "00001111000000000000000000",
        "00011110000000000000000000",
        "00011110000000000000000000",
        "00011110000000000000000000",
        "00011100000000000000000000",
        "00111100001111111100000000",
        "00111101111111111111000000",
        "00111111111111111111100000",
        "00111111111111111111110000",
        "00111111110000000111111000",
        "00111110000000000011111000",
        "00111100000000000001111100",
        "00111100000000000000111100",
        "00111100000000000000111100",
        "00111100000000000000111100",
        "00111100000000000000111100",
        "00111110000000000000111100",
        "00011110000000000000111100",
        "00011110000000000001111000",
        "00011111000000000001111000",
        "00001111100000000011111000",
        "00001111110000001111110000",
        "00000111111111111111100000",
        "00000011111111111111000000",
        "00000001111111111110000000",
        "00000000011111110000000000");
    constant seven: char := (
        "00000000000000000000000000",
        "00111111111111111111111100",
        "00111111111111111111111100",
        "00111111111111111111111100",
        "00111111111111111111111100",
        "00000000000000000001111100",
        "00000000000000000001111000",
        "00000000000000000011111000",
        "00000000000000000011110000",
        "00000000000000000111110000",
        "00000000000000000111100000",
        "00000000000000001111100000",
        "00000000000000001111000000",
        "00000000000000011111000000",
        "00000000000000011111000000",
        "00000000000000111110000000",
        "00000000000000111110000000",
        "00000000000001111100000000",
        "00000000000001111100000000",
        "00000000000011111000000000",
        "00000000000011111000000000",
        "00000000000011110000000000",
        "00000000000111110000000000",
        "00000000000111100000000000",
        "00000000001111100000000000",
        "00000000001111000000000000",
        "00000000011111000000000000",
        "00000000011110000000000000",
        "00000000111110000000000000",
        "00000000111100000000000000",
        "00000001111100000000000000",
        "00000001111100000000000000",
        "00000011111000000000000000",
        "00000011111000000000000000",
        "00000000000000000000000000");
    constant eight: char := (
        "00000000011111111000000000",
        "00000001111111111111000000",
        "00000011111111111111100000",
        "00000111111111111111110000",
        "00001111110000001111110000",
        "00001111000000000011111000",
        "00011110000000000001111000",
        "00011110000000000001111000",
        "00011110000000000001111000",
        "00011110000000000001111000",
        "00011110000000000001111000",
        "00011111000000000011110000",
        "00001111100000000111110000",
        "00000111111000001111100000",
        "00000111111100111111000000",
        "00000011111111111110000000",
        "00000000111111111100000000",
        "00000000111111111100000000",
        "00000001111111111111000000",
        "00000111111100111111100000",
        "00001111110000011111110000",
        "00001111100000000111111000",
        "00011111000000000011111000",
        "00111111000000000011111100",
        "00111110000000000001111100",
        "00111110000000000001111100",
        "00111110000000000001111100",
        "00111110000000000001111100",
        "00111111000000000001111100",
        "00111111000000000011111000",
        "00011111110000001111111000",
        "00001111111111111111110000",
        "00000111111111111111100000",
        "00000011111111111111000000",
        "00000000011111111000000000");
    constant nine: char := (
        "00000000001111111000000000",
        "00000001111111111110000000",
        "00000011111111111111000000",
        "00000111111111111111100000",
        "00001111110000001111110000",
        "00011111000000000111110000",
        "00011110000000000011111000",
        "00011110000000000001111000",
        "00111100000000000001111000",
        "00111100000000000001111000",
        "00111100000000000000111100",
        "00111100000000000000111100",
        "00111100000000000000111100",
        "00111100000000000000111100",
        "00111110000000000000111100",
        "00011111000000000001111100",
        "00011111100000001111111100",
        "00001111111111111111111100",
        "00000111111111111111111100",
        "00000011111111111110111100",
        "00000000111111110000111100",
        "00000000000000000000111000",
        "00000000000000000001111000",
        "00000000000000000001111000",
        "00000000000000000001111000",
        "00000000000000000011110000",
        "00000000000000000111110000",
        "00000000000000001111100000",
        "00000000000000011111000000",
        "00000000000011111111000000",
        "00001111111111111110000000",
        "00001111111111111000000000",
        "00001111111111100000000000",
        "00001111111100000000000000",
        "00000000000000000000000000");
    constant period: char := (
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000111100000000000000000",
        "00001111110000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00001111110000000000000000",
        "00000111100000000000000000");
    constant colon: char := (
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000111100000000000000000",
        "00001111110000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00001111110000000000000000",
        "00000111100000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000000000000000000000000",
        "00000111100000000000000000",
        "00001111110000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00011111111000000000000000",
        "00001111110000000000000000",
        "00000111100000000000000000");
begin
    process(clk, reset) begin
        if (reset = '1') then
            bitline <= (others => '0');
        elsif rising_edge(clk) then
            case bcd is
                when "0000" =>
                    bitline <= zero(to_integer(unsigned(line_num)));
                when "0001" =>
                    bitline <= one(to_integer(unsigned(line_num)));
                when "0010" =>
                    bitline <= two(to_integer(unsigned(line_num)));
                when "0011" =>
                    bitline <= three(to_integer(unsigned(line_num)));
                when "0100" =>
                    bitline <= four(to_integer(unsigned(line_num)));
                when "0101" =>
                    bitline <= five(to_integer(unsigned(line_num)));
                when "0110" =>
                    bitline <= six(to_integer(unsigned(line_num)));
                when "0111" =>
                    bitline <= seven(to_integer(unsigned(line_num)));
                when "1000" =>
                    bitline <= eight(to_integer(unsigned(line_num)));
                when "1001" =>
                    bitline <= nine(to_integer(unsigned(line_num)));
                when "1010" =>
                    bitline <= period(to_integer(unsigned(line_num)));
                when "1011" =>
                    bitline <= colon(to_integer(unsigned(line_num)));
                when others =>
            end case;
        end if;
    end process;
end;
